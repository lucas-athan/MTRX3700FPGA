module hello;
  initial begin
    $display("Hello, Icarus!");
    $finish;
  end
endmodule
